module phase_driver #(
    parameters
) (
    ports
);
    
endmodule